----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    06:05:02 07/28/1963 
-- Design Name: 
-- Module Name:    command_converter - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use ieee.numeric_std.all;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity command_converter is
	Port(command      : in  std_logic_vector(15 downto 0);
		 x             : out std_logic_vector(3  downto 0);
		 y             : out std_logic_vector(3  downto 0);
		 tile          : out std_logic_vector(4  downto 0);
		 piece_bitmap  : out std_logic_vector(24 downto 0));
end command_converter;

architecture Behavioral of command_converter is
	type Matrix is array (0 to 20, 0 to 7) of std_logic_vector(24 downto 0);
	constant piece_lut : Matrix := (
		--a
		 ("0000000000001000000000000",
			"0000000000001000000000000",
			"0000000000001000000000000",
			"0000000000001000000000000",
			"0000000000001000000000000",
			"0000000000001000000000000",
			"0000000000001000000000000",
			"0000000000001000000000000"),
		--b
		("0000000000001000010000000",
			"0000000000001000010000000",
			"0000000000011000000000000",
			"0000000000001100000000000",
			"0000000100001000000000000",
			"0000000100001000000000000",
			"0000000000001100000000000",
			"0000000000011000000000000"),
		--c
		("0000000100001000010000000",
			"0000000100001000010000000",
			"0000000000011100000000000",
			"0000000000011100000000000",
			"0000000100001000010000000",
			"0000000100001000010000000",
			"0000000000011100000000000",
			"0000000000011100000000000"),
		--d
		("0000000100001100000000000",
			"0000000100011000000000000",
			"0000000000001100010000000",
			"0000000000011000010000000",
			"0000000000011000010000000",
			"0000000000001100010000000",
			"0000000100011000000000000",
			"0000000100001100000000000"),
		--e
		("0000000100001000010000100",
			"0000000100001000010000100",
			"0000000000111100000000000",
			"0000000000011110000000000",
			"0100000100001000010000000",
			"0100000100001000010000000",
			"0000000000011110000000000",
			"0000000000111100000000000"),
		--f
		("0000000100001000110000000",
			"0000000100001000011000000",
			"0000001000011100000000000",
			"0000000010011100000000000",
			"0000000110001000010000000",
			"0000001100001000010000000",
			"0000000000011100001000000",
			"0000000000011100100000000"),
		--g
		("0000000100001100010000000",
			"0000000100011000010000000",
			"0000000000011100010000000",
			"0000000000011100010000000",
			"0000000100011000010000000",
			"0000000100001100010000000",
			"0000000100011100000000000",
			"0000000100011100000000000"),
		--h
		("0000000000001100011000000",
			"0000000000011000110000000",
			"0000000000011000110000000",
			"0000000000001100011000000",
			"0000001100011000000000000",
			"0000000110001100000000000",
			"0000000110001100000000000",
			"0000001100011000000000000"),
		--i
		("0000000000011000011000000",
			"0000000000001100110000000",
			"0000000100011000100000000",
			"0000000100001100001000000",
			"0000001100001100000000000",
			"0000000110011000000000000",
			"0000000010001100010000000",
			"0000001000011000010000000"),
		--j
		("0010000100001000010000100",
			"0010000100001000010000100",
			"0000000000111110000000000",
			"0000000000111110000000000",
			"0010000100001000010000100",
			"0010000100001000010000100",
			"0000000000111110000000000",
			"0000000000111110000000000"),
		--k
		("0010000100001000110000000",
			"0010000100001000011000000",
			"0000001000011110000000000",
			"0000000010111100000000000",
			"0000000110001000010000100",
			"0000001100001000010000100",
			"0000000000111100001000000",
			"0000000000011110100000000"),
		--l
		("0010000100011000100000000",
			"0010000100001100001000000",
			"0000001100001110000000000",
			"0000000110111000000000000",
			"0000000010001100010000100",
			"0000001000011000010000100",
			"0000000000111000011000000",
			"0000000000001110110000000"),
		--m
		("0000000100011000110000000",
			"0000000100001100011000000",
			"0000001100011100000000000",
			"0000000110011100000000000",
			"0000000110001100010000000",
			"0000001100011000010000000",
			"0000000000011100011000000",
			"0000000000011100110000000"),
		--n
		("0000001100001000110000000",
			"0000000110001000011000000",
			"0000001010011100000000000",
			"0000001010011100000000000",
			"0000000110001000011000000",
			"0000001100001000110000000",
			"0000000000011100101000000",
			"0000000000011100101000000"),
		--o
		("0000000100001100010000100",
			"0000000100011000010000100",
			"0000000000111100010000000",
			"0000000000011110010000000",
			"0010000100011000010000000",
			"0010000100001100010000000",
			"0000000100011110000000000",
			"0000000100111100000000000"),
		--p
		("0000000100001000111000000",
			"0000000100001000111000000",
			"0000001000011100100000000",
			"0000000010011100001000000",
			"0000001110001000010000000",
			"0000001110001000010000000",
			"0000000010011100001000000",
			"0000001000011100100000000"),
		--q
		("0010000100001110000000000",
			"0010000100111000000000000",
			"0000000000001110010000100",
			"0000000000111000010000100",
			"0000000000111000010000100",
			"0000000000001110010000100",
			"0010000100111000000000000",
			"0010000100001110000000000"),
		--r
		("0000001100001100001000000",
			"0000000110011000100000000",
			"0000000010001100110000000",
			"0000001000011000011000000",
			"0000001000011000011000000",
			"0000000010001100110000000",
			"0000000110011000100000000",
			"0000001100001100001000000"),
		--s
		("0000001000011100001000000",
			"0000000010011100100000000",
			"0000000110001000110000000",
			"0000001100001000011000000",
			"0000001000011100001000000",
			"0000000010011100100000000",
			"0000000110001000110000000",
			"0000001100001000011000000"),
		--t
		("0000001000011100010000000",
			"0000000010011100010000000",
			"0000000110011000010000000",
			"0000001100001100010000000",
			"0000000100011100001000000",
			"0000000100011100100000000",
			"0000000100001100110000000",
			"0000000100011000011000000"),
		--u
		("0000000100011100010000000",
			"0000000100011100010000000",
			"0000000100011100010000000",
			"0000000100011100010000000",
			"0000000100011100010000000",
			"0000000100011100010000000",
			"0000000100011100010000000",
			"0000000100011100010000000"));
begin
	x            <= command(15 downto 12);
	y            <= command(11 downto 8);
	tile         <= command(7 downto 3);
	piece_bitmap <= piece_lut(conv_integer(command(7 downto 3)), conv_integer(command(2 downto 0)));
end Behavioral;

